module complex_butterfly_iter_6_clk_cycles #(
	parameter IWL1 				= 16,
	parameter IWL2 				= 16,
	parameter AWL 				= 17,
	parameter OWL 				= 16,
	parameter CONSTANT_SHIFT	= 1
)(
	input 	wire 				clk,
	input 	wire 				rst,
	input 	wire 				strb_in,
	input 	wire 	[IWL1-1:0]	din1_re,
	input 	wire 	[IWL1-1:0]	din1_im,
	input 	wire 	[IWL2-1:0]	din2_re,
	input 	wire 	[IWL2-1:0]	din2_im,
	input 	wire 	[IWL1-1:0]	din3_re,
	input 	wire 	[IWL1-1:0]	din3_im,
	output 	reg  	[OWL-1:0]	dout1_re,
	output 	reg  	[OWL-1:0]	dout1_im,
	output 	reg  	[OWL-1:0]	dout2_re,
	output 	reg  	[OWL-1:0]	dout2_im,
	output 	wire				strb_out
);
	localparam PROD_WL = IWL1 + IWL2;

	wire	signed	[IWL1-1:0]			MUL_din1_mux;
	wire	signed	[IWL2-1:0]			MUL_din2_mux;

	reg		signed	[PROD_WL-1:0]		tmp_mult;
	reg		signed	[AWL:0]				tmp_mult_out;
	wire			[AWL:0]				mult_out;

	reg				[AWL:0]				mult_reg_1;
	reg				[AWL:0]				mult_reg_2;
	

	wire 			[AWL:0]				pre_sum_din3_re;
	wire 			[AWL:0]				pre_sum_din3_im;

	wire 			[AWL:0]				pre_sum_re_reg;
	wire 			[AWL:0]				pre_sum_im_reg;

	wire	signed	[AWL:0]				ADD_1_din1_mux;
	wire	signed	[AWL:0]				ADD_1_din2_mux;

	wire	signed	[AWL:0]				SUB_1_din1_mux; 
	wire	signed	[AWL:0]				SUB_1_din2_mux;

	reg		signed	[AWL:0]				tmp_add_1;
	reg		signed	[AWL:0]				tmp_sub_1;

	reg				[OWL-1:0]			add_1_out;
	reg				[OWL-1:0]			sub_1_out;

	reg				[OWL-1:0]			re_reg;
	reg				[OWL-1:0]			im_reg;

	reg			  	[OWL-1:0]			dout1_re_b;
	reg			  	[OWL-1:0]			dout2_re_b;

	reg				[2:0]				pipe_cnt;
	wire								valid;

	assign valid 		= 	pipe_cnt[2] && pipe_cnt[0];

	assign strb_out		= 	strb_in;


	always @(posedge clk) begin : pipe_alw
		if(rst) begin
			pipe_cnt <= 0;
		end else begin 
			if(strb_in) begin 
				pipe_cnt <= 0;
			end else begin
				if (!(pipe_cnt[2] && pipe_cnt[0])) begin
					pipe_cnt <= pipe_cnt + 1;
				end
			end
		end
	end

	assign MUL_din1_mux	=	(pipe_cnt[0])				? 	din1_im	: din1_re;
	assign MUL_din2_mux	=	(pipe_cnt[0] ^ pipe_cnt[1])	? 	din2_im	: din2_re;

	always @(*) begin : mult_alw
		tmp_mult = MUL_din1_mux * MUL_din2_mux;
		tmp_mult_out = tmp_mult[PROD_WL-1:PROD_WL-AWL-1];
	end

	assign mult_out 		= (CONSTANT_SHIFT == 0)? tmp_mult_out :  tmp_mult_out >>> 1;
	
	assign pre_sum_din3_re 	= (CONSTANT_SHIFT == 0)? {din3_re[IWL1-1], din3_re, 1'b0}: {din3_re[IWL1-1], din3_re[IWL1-1], din3_re};
	assign pre_sum_din3_im 	= (CONSTANT_SHIFT == 0)? {din3_im[IWL1-1], din3_im, 1'b0}: {din3_im[IWL1-1], din3_im[IWL1-1], din3_im};
	
	assign pre_sum_re_reg 	= {re_reg[OWL-1], re_reg, 1'b0};
	assign pre_sum_im_reg 	= {im_reg[OWL-1], im_reg, 1'b0};

	assign ADD_1_din1_mux =	(pipe_cnt[2])? 	((pipe_cnt[0])? pre_sum_im_reg : mult_reg_1)	:	pre_sum_re_reg ;
	assign ADD_1_din2_mux =	(pipe_cnt[2])? 	((pipe_cnt[0])? pre_sum_din3_im : mult_reg_2)	:	pre_sum_din3_re ;


	always @* begin : add_1_alw
		tmp_add_1 = ADD_1_din1_mux + ADD_1_din2_mux + 2'b01;
		if (tmp_add_1[AWL] == tmp_add_1[AWL-1]) begin 
			add_1_out = tmp_add_1[AWL-1: AWL-OWL];
		end else begin 
			add_1_out[OWL-1] = tmp_add_1[AWL];
			add_1_out[OWL-2:0] = {OWL-1{tmp_add_1[AWL-1]}};
		end 
	end

	assign SUB_1_din2_mux =	(pipe_cnt[2])? pre_sum_im_reg 	: ((pipe_cnt[0])? pre_sum_re_reg : mult_reg_1);
	assign SUB_1_din1_mux =	(pipe_cnt[2])? pre_sum_din3_im	: ((pipe_cnt[0])? pre_sum_din3_re : mult_reg_2);


	always @* begin : sub_1_alw
		tmp_sub_1 = SUB_1_din1_mux - SUB_1_din2_mux + 2'b01;
		if (tmp_sub_1[AWL] == tmp_sub_1[AWL-1]) begin 
			sub_1_out = tmp_sub_1[AWL-1: AWL-OWL];
		end else begin 
			sub_1_out[OWL-1] = tmp_sub_1[AWL];
			sub_1_out[OWL-2:0] = {OWL-1{tmp_sub_1[AWL-1]}};
		end 
	end


	
	always @(posedge clk) begin : pipe_mult_reg1
		if(!(pipe_cnt[0] | pipe_cnt[2])) begin 
			mult_reg_1 <= mult_out;
		end
	end

	always @(posedge clk) begin : pipe_mult_reg2
		if(pipe_cnt[0] & ~pipe_cnt[2]) begin 
			mult_reg_2 <= mult_out;
		end
	end

	always @(posedge clk) begin
		if(pipe_cnt == 3'b010) begin 
			re_reg <= sub_1_out;
		end
	end

	always @(posedge clk) begin
		if(pipe_cnt == 3'b100) begin 
			im_reg <= add_1_out;
		end
	end

	always @(posedge clk) begin
		if(pipe_cnt == 3'b011) begin 
			dout1_re_b <= add_1_out; 
			dout2_re_b <= sub_1_out;
		end
	end


	always @(posedge clk) begin
		if(rst) begin
			dout1_re <= 0;
			dout1_im <= 0;
			dout2_re <= 0;
			dout2_im <= 0;
		end else begin 
			if(strb_in && valid) begin
				dout2_re <= dout1_re_b;
				dout1_im <= add_1_out;
				dout1_re <= dout2_re_b;
				dout2_im <= sub_1_out;
			end
		end
	end


endmodule 		
			
	